module accelerator_tb();


endmodule
